* SPICE NETLIST
***************************************

.SUBCKT XOR2 GND VDD I[1] I[2] I[3] I[4] out
** N=10 EP=7 IP=0 FDC=8
* PORT GND GND 30000 2500 METAL3
* PORT VDD VDD 30000 57500 METAL3
* PORT I[1] I[1] 12500 31000 METAL3
* PORT I[2] I[2] 23500 31000 METAL3
* PORT I[3] I[3] 35000 30500 METAL3
* PORT I[4] I[4] 49000 23000 METAL3
* PORT out out 57500 30000 METAL3
M0 9 I[1] GND GND N L=1.8e-07 W=5.4e-07 AD=1.944e-13 AS=2.5515e-13 $X=19000 $Y=11000 $D=1
M1 out I[2] 9 GND N L=1.8e-07 W=5.4e-07 AD=2.916e-13 AS=1.944e-13 $X=25000 $Y=11000 $D=1
M2 10 I[3] out GND N L=1.8e-07 W=5.4e-07 AD=1.944e-13 AS=2.916e-13 $X=33000 $Y=11000 $D=1
M3 GND I[4] 10 GND N L=1.8e-07 W=5.4e-07 AD=2.5515e-13 AS=1.944e-13 $X=39000 $Y=11000 $D=1
M4 8 I[1] VDD VDD P L=1.8e-07 W=1.08e-06 AD=5.832e-13 AS=5.2245e-13 $X=13000 $Y=36000 $D=0
M5 VDD I[2] 8 VDD P L=1.8e-07 W=1.08e-06 AD=5.2245e-13 AS=5.832e-13 $X=21000 $Y=36000 $D=0
M6 out I[3] 8 VDD P L=1.8e-07 W=1.08e-06 AD=5.832e-13 AS=5.346e-13 $X=37000 $Y=36000 $D=0
M7 8 I[4] out VDD P L=1.8e-07 W=1.08e-06 AD=6.318e-13 AS=5.832e-13 $X=45000 $Y=36000 $D=0
.ENDS
***************************************
